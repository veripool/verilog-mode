// msg1354
module f (/*AUTOARG*/
          // Outputs
          o2,
          o1,
          // Inputs
          z,
          a,
          q
          );
   
   output o2;
   input  z;
   input  a;
   input  q;
   output o1;
endmodule

// Local Variables:
// verilog-auto-arg-format:single
// End:
