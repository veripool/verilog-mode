module mymodule();
   parameter real fc=10e6;
   parameter real bw=25e3;
   
   analog begin
      // contents of module here
   end // analog
   
endmodule // mymodule

// Local Variables:
// verilog-minimum-comment-distance: 1
// verilog-auto-endcomments: t
// End:
