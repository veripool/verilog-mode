module autoinoutin (/*AUTOARG*/
                    // Inputs
                    lower_inb, lower_ina, lower_out
                    );
   
   /*AUTOINOUTIN("inst")*/
   // Beginning of automatic in/out/inouts (from specific module)
   input lower_inb;
   input lower_ina;
   input lower_out;
   // End of automatics
   
endmodule

