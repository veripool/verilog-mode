module top
  (
   /*AUTOOUTPUTEVERY("^a")*/
   // Beginning of automatic outputs (every signal)
   output aa,
   output ab
   // End of automatics
   );
   
   wire aa;
   wire ab;
   wire cc;
endmodule
