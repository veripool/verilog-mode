module ocnSwitchClockGen(output reg ocnSwitchClock);
   parameter   ocnSwitchClockPeriod = 2000;
