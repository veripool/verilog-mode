parameter
  // full line comment
  param1 = 1'b1,  // trailing comment
  param2 = 1'b0,  /* trailing comment */
         // full line comment
  param3 = 1'b1;
