module tahoetop(/*AUTOARG*/);

   /*AUTOWIRE*/
   // Beginning of automatic wires (for undeclared instantiated-module outputs)
   // End of automatics


   // the pad instance to look like "pads pads (/*AUTOINST*/". Then at
   // diff the new against the old. Finally delete /*AUTOINST*/. This will

endmodule
