module foo # (
parameter A = 0,
parameter B = 0,
parameter C = 0,
parameter D = 0
)(
input wire a,
input wire b,
output reg z
);
endmodule


// Local Variables:
// verilog-indent-lists: nil
// End:
