module ex;

   /* autoinst_paramover_sub AUTO_TEMPLATE "u_\(.*\)" (
    .a(inA_@[]),
    .b(outA_@[]),
    );*/

   autoinst_paramover_sub u_foo(/*AUTOINST*/);
   autoinst_paramover_sub u_bar(/*AUTOINST*/);
   autoinst_paramover_sub u_baz(/*AUTOINST*/);

   /* autoinst_paramover_sub AUTO_TEMPLATE (
    .a(inN_@[]),
    .b(outN_@[]),
    );*/

   autoinst_paramover_sub u_0_2(/*AUTOINST*/);
   autoinst_paramover_sub u_1_3(/*AUTOINST*/);

endmodule
