module ExampArg (/*AUTOARG*/
                 // Outputs
                 o,
                 // Inputs
                 i
                 );
   input  i;
   output o;
endmodule

// Local Variables:
// indent-tabs-mode: nil
// End:
