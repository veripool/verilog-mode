module ExampInsertLisp;

   /*AUTOINSERTLAST(my-verilog-insert-hello "world")*/

endmodule
/*
 Local Variables:
 eval:
   (defun my-verilog-insert-hello (who)
     (insert (concat "initial $write(\"hello " who "\");\n")))
 End:
*/
