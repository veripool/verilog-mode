module foo(reg_input_signal_name,a,b,c,d,e);
   // foo bar
   output 	     c;//this is a comment


   reg 		     foo;
   //a

   /*  jj
    KK */
   reg 		     foo;
   output        reg /*   */  signed 	     d;
   output reg signed e; /* so is this */

   reg [31:0] 	     blather;

endmodule // foo

