module top
  (
   /*AUTOOUTPUTEVERY("^a")*/
   );   

   wire 		aa;
   wire 		ab;
   wire 		cc;
endmodule
