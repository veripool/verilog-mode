module Ptest #(
       parameter I_CONTROL     = 8'h 00, R_CONTROL     = 8'h00)
  ( 
   input scanTest,
   input scanArst);
endmodule 

module t;

  Ptest
    #(/*AUTOINSTPARAM*/)
   u_Ptest
     (/*AUTOINST*/);

endmodule
