module autoinoutmodule_iface_sub
  (my_svi.master my_svi_port,
   );
endmodule
