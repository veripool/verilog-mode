module autowire_topv_two;
   output logic [1:0] foo2;
endmodule
