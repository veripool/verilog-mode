module autoinoutmodule_re2 (/*AUTOARG*/);

   /*AUTOINOUTMODULE("inst","","input.*")*/

   /*AUTOINOUTMODULE("inst","","output.*")*/

   wire   lower_out  = lower_ina;

endmodule

