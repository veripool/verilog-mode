
module flag_f_reeves
  (/*AUTOARG*/) ;

   /*AUTOOUTPUT*/

   /*AUTOINPUT*/

   flag_f_reeves_IBUF ibuf
     (/*AUTOINST*/);

endmodule
// Local Variables:
// verilog-library-flags: ("-f flag_f_reeves.vc")
// End:
