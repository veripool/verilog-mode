module autowire_topv_one;
   output [1:0] foo;
   output [1:0] bar;
endmodule
