module lavigne_t2 (b);
input b;
endmodule
