module batch_prof_cell(Z,A,B);
   output Z;
   input  A, B;
endmodule
