module aaa();
   always @(a) begin
      if (a) begin
         /*AUTORESET*/
      end
      // note missing e-n-d
   always @(*) begin
   end
endmodule
