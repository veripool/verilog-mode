        module ExampArg (/*AUTOARG*/);
          input i;
          output o;
        endmodule

// Local Variables:
// indent-tabs-mode: nil
// End:
