module autowire_long_yaohung(/*AUTOARG*/);
   
   /*AUTOOUTPUT*/
   /*AUTOWIRE*/
   /*AUTOREG*/
   
   top top
     (/*AUTOINST*/);
   
endmodule

module top(/*AUTOARG*/);
   
   output [`LONGNAMELONGNAMELONGNAMELONGNAMELONGNAMELONGNAME] data_out;
   
endmodule
