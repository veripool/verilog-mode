module autoinoutmodule (/*AUTOARG*/);

   /*AUTOINOUTMODULE("inst","ina\|out")*/
   // Beginning of automatic in/out/inouts (from specific module)

   wire   lower_out = lower_ina;

endmodule

