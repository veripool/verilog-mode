input  bar;
output foo;
