module (/*AUTOARG*/
        // Outputs
        o1, o2,
        // Inputs
        a, q, z
        );
   output o2;
   input  z;
   input  a;
   input  q;
   output o1;
endmodule

// Local Variables:
// verilog-auto-arg-sort:t
// End:
