module autowire_topv_two;
   output logic [1:0] foo2;
   output logic       foo3;
   output logic [1:0] bar2;
   output logic       bar3;
endmodule
