// bug360
module f (/*AUTOARG*/
          // Inputs
          x
          );
   
   always @* r = "test/*";
   
   input x;
   
endmodule
