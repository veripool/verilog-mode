module autoinoutmodule (/*AUTOARG*/);

   /*AUTOINOUTMODULE("inst","ina\|out")*/

   wire   lower_out = lower_ina;

endmodule

