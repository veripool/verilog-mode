// bug360
module f (/*AUTOARG*/);

always @* r = "test/*";

  input 				x;

endmodule
