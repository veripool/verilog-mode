`include "some_macros.v"

module z();
  
   $display("%t:", $time);
   a 			      = b;
   casfasdf 		      = d;
   g 			      = r;
   fgasdfasdfasdfasfdasfd    <= p;
   gh 			     := h;
   gf 			     <=g;
   ssdf 		      = 5;
   f 			      = zsfdsdf >= f;
  
endmodule
