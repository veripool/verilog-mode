module tahoetop(/*AUTOARG*/);
   
   /*AUTOWIRE*/
   
   
   // the pad instance to look like "pads pads (/*AUTOINST*/". Then at
   // diff the new against the old. Finally delete /*AUTOINST*/. This will
   
endmodule
