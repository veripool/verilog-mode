module lavigne_t1 (a);
input a;
endmodule
