// bug 841
module x;

always @*
begin
end // always @ *

endmodule // x

// Local Variables:
// verilog-indent-level-module: 0
// verilog-indent-begin-after-if: nil
// verilog-minimum-comment-distance: 1
// verilog-auto-endcomments: t
// End:
