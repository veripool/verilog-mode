// bug721
module my_core
  (
   /*AUTOINOUTMODULE("autoinoutmodule_iface_sub")*/
   /*AUTOINOUT*/
   /*AUTOINPUT*/
   /*AUTOOUTPUT*/
);
/*AUTOWIRE*/

endmodule
