module x;
   parameter Pp = 1;
   /*AUTOINSERTLISP(insert vh-Pp "\n")*/
   // Beginning of automatic insert lisp
   1
     // End of automatics
     
     localparam Lp = 2;
   /*AUTOINSERTLISP(insert vh-Lp "\n")*/
   // Beginning of automatic insert lisp
   2
     // End of automatics
     
     parameter mytype_t Pt = 3;
   /*AUTOINSERTLISP(insert vh-Pt "\n")*/
   // Beginning of automatic insert lisp
   3
     // End of automatics
     
     endmodule

// Local Variables:
// verilog-library-directories: (".")
// eval:(verilog-read-defines)
// End:
