module x;
   parameter Pp = 1;
   /*AUTOINSERTLISP(insert vh-Pp "\n")*/

   localparam Lp = 2;
   /*AUTOINSERTLISP(insert vh-Lp "\n")*/

   parameter mytype_t Pt = 3;
   /*AUTOINSERTLISP(insert vh-Pt "\n")*/

endmodule

// Local Variables:
// verilog-library-directories: (".")
// eval:(verilog-read-defines)
// End:
