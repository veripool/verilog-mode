module autoinstparam_belkind_leaf (/*AUTOARG*/
   // Inputs
   a
   ) ;

   parameter P =3D 4;
   input [P-1:0] a;

endmodule // leaf
// Local Variables:
// eval:(verilog-read-defines)
// End:
