module autoinst_ifdef_fredrickson_200503_top();

   autoinst_ifdef_fredrickson_200503_sub sub
    (/*AUTOINST*/
     // Outputs
     .d					(d),
     .b					(b),
     // Inputs
     .a					(a),
     .c					(c));

endmodule // define_top
