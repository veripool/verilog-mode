module autowire_topv;
   /*AUTOOUTPUT("bar")*/

   /*AUTOWIRE*/

   autowire_topv_one one (/*AUTOINST*/);
   autowire_topv_two two (/*AUTOINST*/);
endmodule

// Local Variables:
// verilog-auto-wire-type: "wire"
// End:
