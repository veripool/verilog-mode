module autoinstparam_belkind_leaf (/*AUTOARG*/) ;

   parameter P =3D 4;
   input [P-1:0] a;

endmodule // leaf
// Local Variables:
// verilog-auto-read-includes:t
// End:
