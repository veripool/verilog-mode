module autoinoutparam (/*AUTOARG*/);

   /*AUTOINOUTPARAM("inst","param1")*/

   /*AUTOINOUTPARAM("inst")*/

endmodule

