// bug721
module my_core
  (
   /*AUTOINOUTMODULE("autoinoutmodule_iface_sub")*/
   // Beginning of automatic in/out/inouts (from specific module)
   my_svi.master my_svi_port
   // End of automatics
   /*AUTOINOUT*/
   /*AUTOINPUT*/
   /*AUTOOUTPUT*/
   );
   /*AUTOWIRE*/
   
endmodule
