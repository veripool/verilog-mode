// bug 842
module x;

do begin
end while();

endmodule

// Local Variables:
// verilog-minimum-comment-distance: 1
// verilog-auto-endcomments: t
// End:
