module autoinoutmodule (
   /*AUTOINOUTMODULE("inst")*/
   );

   wire   lower_out = lower_ina | lower_inb;

endmodule

