module autoinst_sv_shaw
  (
   /*AUTOINOUTMODULE("Example_mod")*/
   );

   Example_mod Ex1 (/*AUTOINST*/);

endmodule

module Example_mod
  (
    input  logic clk,
    input  logic reset_b,
   );
endmodule

