module io1_sub(
   /*AUTOINPUT*/
   /*AUTOOUTPUT*/
   );

   /* inst AUTO_TEMPLATE (
    .lower_inb		(1'b1),
    )*/


   inst inst (/*AUTOINST*/);

endmodule
