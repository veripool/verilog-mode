module top;
   /*AUTOWIRE*/
   sub0 #(/*AUTOINSTPARAM*/)
   s0 (/*AUTOINST*/);
endmodule

module sub0
  #(
    parameter string testit2 = 0,
    int TESTIT = 0
    ) (
       // clk and resets
    input  logic   side_clk,
    input  logic   side_rst_b,
       );

endmodule
