package p;
typedef enum {a, b} type_t;
typedef enum {TASK, TASK2} type2_t;
typedef enum {Package, Class} type3_t;
endpackage
