// bug 825
module x;

always @*
begin
end

initial
begin
end

final
begin
end

endmodule

// Local Variables:
// verilog-indent-begin-after-if: nil
// End:
