module foo # (
   parameter A = 0,
   B           = 0,
   C           = 0,
   D           = 0
)(
   input wire a,
   input wire b,
   output reg z
);
endmodule


// Local Variables:
// verilog-indent-lists: nil
// End:
