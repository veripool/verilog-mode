module autoinoutparam (/*AUTOARG*/);
   
   /*AUTOINOUTPARAM("inst","param1")*/
   // Beginning of automatic parameters (from specific module)
   parameter param1;
   // End of automatics
   
   /*AUTOINOUTPARAM("inst")*/
   // Beginning of automatic parameters (from specific module)
   parameter param2;
   // End of automatics
   
endmodule

