// msg1354
module f (/*AUTOARG*/);

   output o2;
   input z;
   input a;
   input q;
   output o1;
endmodule

// Local Variables:
// verilog-auto-arg-format:single
// End:
