// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2011 by Wilson Snyder.

// Note intentional whitespace on following line
//       SPACES
module x;      
   //       TAB
endmodule	

// Local Variables:
// verilog-auto-delete-trailing-whitespace: t
// End:
