module top
  (
   /*AUTOINPUT*/
   );

   /*AUTOWIRE*/

   inst_module inst (/*AUTOINST*/);
endmodule

module inst_module (input supply0 VDD,
                    input supply1 VSS,
		    input non_supply,
		    input supply1 VDD_from_child
		    );

endmodule
