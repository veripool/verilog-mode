module autoinoutmodule (/*AUTOARG*/);

   /*AUTOINOUTMODULE("inst","\(ina\|out\)","","ina")*/

   wire   lower_out = lower_ina;

endmodule

