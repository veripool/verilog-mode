interface class ic;
   // ...
endclass
// this should indent to left margin, but indented one stop to right
