module (/*AUTOARG*/);
   output o2;
   input z;
   input a;
   input q;
   output o1;
endmodule

// Local Variables:
// verilog-auto-arg-sort:t
// End:
