// Bug 888 -- verilog-label-be should remove existing comment labels before adding new ones
class c;
endclass // delete-me
