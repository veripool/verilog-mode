module TEST_TOP (
                 );
   /*TEST AUTO_TEMPLATE
    (
    
    .abcd_efgh_ijklmno_f02_out_c(abcdefg_f02_clroilouull[5]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_be_2(abcdefg_f10_eg2_ab_cdefghijklm[49]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_fh_2(abcdefg_f08_eg0_ab_a_fghi[6]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_ch(abcdefg_f09_eg1_ab_cdefghijklm[36]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_ej_1(abcdefg_f10_eg2_ab_cdefghijklm[14]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_ga_1(abcdefg_f10_eg2_ab_cdefghijklm[3]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_fe(abcdefg_f09_eg1_ab_cdefghijklm[9]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_bi_2(abcdefg_f08_eg0_ab_cdefghijklm[45]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_24_1(abcdefg_f09_eg1_ab_fghijklm[24]),
    .abcd_efgh_ijklmno_f01_oilouull_o_0_1(abcdefg_f01_oilouull[0]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_cc_2(abcdefg_f10_eg2_ab_cdefghijklm[41]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_e_2(abcdefg_f11_eg3_ab_cdefghijklm[59]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_54_1(abcdefg_f11_eg3_ab_fghijklm[54]),
    .abcd_efgh_ijklmno_f03_oilouull_o_3_1(abcdefg_f03_oilouull[3]),
    .abcd_efgh_ijklmno_f02_out_h_2(abcdefg_f02_a_zxdf[0]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_g_1(abcdefg_f11_eg3_ab_a_fghi[57]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_b_2(abcdefg_f08_eg0_ab_cdefghijklm[62]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_9_1(abcdefg_f11_eg3_ab_fghijklm[9]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_di_1(abcdefg_f09_eg1_ab_a_fghi[25]),
    .abcd_efgh_ijklmno_f00_out_h_2(abcdefg_f00_a_zxdf[0]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_cg_2(abcdefg_f11_eg3_ab_cdefghijklm[37]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_eh_2(abcdefg_f10_eg2_ab_a_fghi[16]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_di_1(abcdefg_f08_eg0_ab_cdefghijklm[25]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_ec_2(abcdefg_f11_eg3_ab_cdefghijklm[21]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_d_1(abcdefg_f11_eg3_ab_a_fghi[60]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_bh_1(abcdefg_f11_eg3_ab_a_fghi[46]),
    .abcd_efgh_ijklmno_f00_out_f(abcdefg_f00_clroilouull[2]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_52_1(abcdefg_f11_eg3_ab_fghijklm[52]),
    .abcd_efgh_ijklmno_f02_out_g(abcdefg_f02_clroilouull[1]),
    .abcd_efgh_ijklmno_f07_out_e(abcdefg_f07_clroilouull[3]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_ff_2(abcdefg_f10_eg2_ab_a_fghi[8]),
    .abcd_efgh_ijklmno_f04_out_h(abcdefg_f04_clroilouull[0]),
    .abcd_efgh_ijklmno_f04_out_g_2(abcdefg_f04_a_zxdf[1]),
    .abcd_efgh_ijklmno_f02_out_c_2(abcdefg_f02_a_zxdf[5]),
    .abcd_efgh_ijklmno_f04_out_a_3(abcdefg_f04_a_zxdf[7]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_fa_1(abcdefg_f08_eg0_ab_cdefghijklm[13]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_ed_2(abcdefg_f08_eg0_ab_a_fghi[20]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_ea_2(abcdefg_f10_eg2_ab_a_fghi[23]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_c_2(abcdefg_f10_eg2_ab_cdefghijklm[61]),
    .abcd_efgh_ijklmno_f03_oilouull_o_0_1(abcdefg_f03_oilouull[0]),
    .abcd_efgh_ijklmno_f00_out_e_2(abcdefg_f00_a_zxdf[3]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_bg_3(abcdefg_f10_eg2_ab_a_fghi[47]),
    .abcd_efgh_ijklmno_f05_oilouull_o_2_1(abcdefg_f05_oilouull[2]),
    .abcd_efgh_ijklmno_f01_out_h_2(abcdefg_f01_a_zxdf[0]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_44_1(abcdefg_f10_eg2_ab_fghijklm[44]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_j_3(abcdefg_f08_eg0_ab_a_fghi[54]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_39_1(abcdefg_f08_eg0_ab_fghijklm[39]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_fj_2(abcdefg_f08_eg0_ab_a_fghi[4]),
    .abcd_efgh_ijklmno_f05_out_h(abcdefg_f05_clroilouull[0]),
    .abcd_efgh_ijklmno_f05_out_d_2(abcdefg_f05_a_zxdf[4]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_gb_2(abcdefg_f10_eg2_ab_a_fghi[2]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_cb_3(abcdefg_f10_eg2_ab_a_fghi[42]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_52_1(abcdefg_f10_eg2_ab_fghijklm[52]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_be_2(abcdefg_f11_eg3_ab_cdefghijklm[49]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_42_1(abcdefg_f11_eg3_ab_fghijklm[42]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_ci_1(abcdefg_f11_eg3_ab_a_fghi[35]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_fh_1(abcdefg_f10_eg2_ab_cdefghijklm[6]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_24_1(abcdefg_f08_eg0_ab_fghijklm[24]),
    .abcd_efgh_ijklmno_f02_out_g_2(abcdefg_f02_a_zxdf[1]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_d_2(abcdefg_f11_eg3_ab_cdefghijklm[60]),
    .abcd_efgh_ijklmno_f06_out_d_2(abcdefg_f06_a_zxdf[4]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_ea_1(abcdefg_f09_eg1_ab_a_fghi[23]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_dh_2(abcdefg_f11_eg3_ab_cdefghijklm[26]),
    .abcd_efgh_ijklmno_f04_oilouull_o_7_2(abcdefg_f04_oilouull[7]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_dh_1(abcdefg_f09_eg1_ab_a_fghi[26]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_18_1(abcdefg_f08_eg0_ab_fghijklm[18]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_ba_2(abcdefg_f11_eg3_ab_cdefghijklm[53]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_ce_1(abcdefg_f11_eg3_ab_a_fghi[39]),
    .abcd_efgh_ijklmno_f03_oilouull_o_5_1(abcdefg_f03_oilouull[5]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_ef_1(abcdefg_f09_eg1_ab_a_fghi[18]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_cj_2(abcdefg_f08_eg0_ab_cdefghijklm[34]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_j_2(abcdefg_f08_eg0_ab_cdefghijklm[54]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_bh_3(abcdefg_f08_eg0_ab_a_fghi[46]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_cb_1(abcdefg_f09_eg1_ab_a_fghi[42]),
    .abcd_efgh_ijklmno_f01_oilouull_o_6_2(abcdefg_f01_oilouull[6]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_ba_3(abcdefg_f10_eg2_ab_a_fghi[53]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_0_1(abcdefg_f11_eg3_ab_fghijklm[0]),
    .abcd_efgh_ijklmno_f06_out_h_2(abcdefg_f06_a_zxdf[0]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_51_1(abcdefg_f08_eg0_ab_fghijklm[51]),
    .abcd_efgh_ijklmno_f06_oilouull_o_4_1(abcdefg_f06_oilouull[4]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_10_1(abcdefg_f08_eg0_ab_fghijklm[10]),
    .abcd_efgh_ijklmno_f01_oilouull_o_7_2(abcdefg_f01_oilouull[7]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_da_2(abcdefg_f11_eg3_ab_cdefghijklm[33]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_e_1(abcdefg_f09_eg1_ab_a_fghi[59]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_22_1(abcdefg_f08_eg0_ab_fghijklm[22]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_db_2(abcdefg_f11_eg3_ab_cdefghijklm[32]),
    .abcd_efgh_ijklmno_f01_oilouull_o_2_1(abcdefg_f01_oilouull[2]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_ci_3(abcdefg_f08_eg0_ab_a_fghi[35]),
    .abcd_efgh_ijklmno_f07_oilouull_o_6_2(abcdefg_f07_oilouull[6]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_62_1(abcdefg_f11_eg3_ab_fghijklm[62]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_34_1(abcdefg_f10_eg2_ab_fghijklm[34]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_9_1(abcdefg_f10_eg2_ab_fghijklm[9]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_13_1(abcdefg_f10_eg2_ab_fghijklm[13]),
    .abcd_efgh_ijklmno_f05_oilouull_o_7_2(abcdefg_f05_oilouull[7]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_ch_1(abcdefg_f11_eg3_ab_a_fghi[36]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_fd_1(abcdefg_f10_eg2_ab_cdefghijklm[10]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_fc_2(abcdefg_f10_eg2_ab_a_fghi[11]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_ei_1(abcdefg_f09_eg1_ab_a_fghi[15]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_37_1(abcdefg_f08_eg0_ab_fghijklm[37]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_gb(abcdefg_f09_eg1_ab_cdefghijklm[2]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_7_1(abcdefg_f10_eg2_ab_fghijklm[7]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_dg_2(abcdefg_f11_eg3_ab_cdefghijklm[27]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_ce(abcdefg_f09_eg1_ab_cdefghijklm[39]),
    .abcd_efgh_ijklmno_f07_out_d_2(abcdefg_f07_a_zxdf[4]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_cd_2(abcdefg_f08_eg0_ab_cdefghijklm[40]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_57_1(abcdefg_f10_eg2_ab_fghijklm[57]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_63_1(abcdefg_f10_eg2_ab_fghijklm[63]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_j_1(abcdefg_f09_eg1_ab_a_fghi[54]),
    .abcd_efgh_ijklmno_f00_out_a(abcdefg_f00_clroilouull[7]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_46_1(abcdefg_f09_eg1_ab_fghijklm[46]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_39_1(abcdefg_f10_eg2_ab_fghijklm[39]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_28_1(abcdefg_f08_eg0_ab_fghijklm[28]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_20_1(abcdefg_f08_eg0_ab_fghijklm[20]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_51_1(abcdefg_f11_eg3_ab_fghijklm[51]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_ci_1(abcdefg_f09_eg1_ab_a_fghi[35]),
    .abcd_efgh_ijklmno_f04_out_h_2(abcdefg_f04_a_zxdf[0]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_bd(abcdefg_f09_eg1_ab_cdefghijklm[50]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_dg_1(abcdefg_f10_eg2_ab_cdefghijklm[27]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_23_1(abcdefg_f09_eg1_ab_fghijklm[23]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_1_2(abcdefg_f09_eg1_ab_fghijklm[1]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_bc_2(abcdefg_f08_eg0_ab_cdefghijklm[51]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_bc_3(abcdefg_f10_eg2_ab_a_fghi[51]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_62_1(abcdefg_f08_eg0_ab_fghijklm[62]),
    .abcd_efgh_ijklmno_f01_out_g_2(abcdefg_f01_a_zxdf[1]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_23_1(abcdefg_f11_eg3_ab_fghijklm[23]),
    .abcd_efgh_ijklmno_f03_out_e_2(abcdefg_f03_a_zxdf[3]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_b_1(abcdefg_f09_eg1_ab_a_fghi[62]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_eh(abcdefg_f09_eg1_ab_cdefghijklm[16]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_dh_1(abcdefg_f10_eg2_ab_cdefghijklm[26]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_34_1(abcdefg_f09_eg1_ab_fghijklm[34]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_gc_1(abcdefg_f10_eg2_ab_cdefghijklm[1]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_cg_2(abcdefg_f08_eg0_ab_cdefghijklm[37]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_13_1(abcdefg_f11_eg3_ab_fghijklm[13]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_2_1(abcdefg_f08_eg0_ab_fghijklm[2]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_fb(abcdefg_f09_eg1_ab_cdefghijklm[12]),
    .abcd_efgh_ijklmno_f00_oilouull_o_6_2(abcdefg_f00_oilouull[6]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_h_3(abcdefg_f08_eg0_ab_a_fghi[56]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_38_1(abcdefg_f09_eg1_ab_fghijklm[38]),
    .abcd_efgh_ijklmno_f00_out_c(abcdefg_f00_clroilouull[5]),
    .abcd_efgh_ijklmno_f06_out_a_3(abcdefg_f06_a_zxdf[7]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_60_1(abcdefg_f09_eg1_ab_fghijklm[60]),
    .abcd_efgh_ijklmno_f06_oilouull_o_2_1(abcdefg_f06_oilouull[2]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_8_1(abcdefg_f09_eg1_ab_fghijklm[8]),
    .abcd_efgh_ijklmno_f03_out_f(abcdefg_f03_clroilouull[2]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_dj_1(abcdefg_f08_eg0_ab_cdefghijklm[24]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_bg_2(abcdefg_f08_eg0_ab_cdefghijklm[47]),
    .abcd_efgh_ijklmno_f01_oilouull_o_4_1(abcdefg_f01_oilouull[4]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_ef_2(abcdefg_f10_eg2_ab_a_fghi[18]),
    .abcd_efgh_ijklmno_f01_out_a_3(abcdefg_f01_a_zxdf[7]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_12_1(abcdefg_f08_eg0_ab_fghijklm[12]),
    .abcd_efgh_ijklmno_f07_out_c_2(abcdefg_f07_a_zxdf[5]),
    .abcd_efgh_ijklmno_f00_out_e(abcdefg_f00_clroilouull[3]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_ca_1(abcdefg_f09_eg1_ab_a_fghi[43]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_eg_2(abcdefg_f08_eg0_ab_a_fghi[17]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_be_1(abcdefg_f11_eg3_ab_a_fghi[49]),
    .abcd_efgh_ijklmno_f06_out_d(abcdefg_f06_clroilouull[4]),
    .abcd_efgh_ijklmno_f00_out_g(abcdefg_f00_clroilouull[1]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_b(abcdefg_f09_eg1_ab_cdefghijklm[62]),
    .abcd_efgh_ijklmno_f00_out_f_2(abcdefg_f00_a_zxdf[2]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_gc_1(abcdefg_f09_eg1_ab_a_fghi[1]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_ca_1(abcdefg_f11_eg3_ab_a_fghi[43]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_ea(abcdefg_f09_eg1_ab_cdefghijklm[23]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_12_1(abcdefg_f10_eg2_ab_fghijklm[12]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_gd_2(abcdefg_f11_eg3_ab_cdefghijklm[0]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_i_1(abcdefg_f09_eg1_ab_a_fghi[55]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_e_2(abcdefg_f08_eg0_ab_cdefghijklm[59]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_ff(abcdefg_f09_eg1_ab_cdefghijklm[8]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_17_1(abcdefg_f11_eg3_ab_fghijklm[17]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_be_3(abcdefg_f10_eg2_ab_a_fghi[49]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_20_1(abcdefg_f11_eg3_ab_fghijklm[20]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_bc_1(abcdefg_f11_eg3_ab_a_fghi[51]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_43_1(abcdefg_f09_eg1_ab_fghijklm[43]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_54_1(abcdefg_f09_eg1_ab_fghijklm[54]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_be_2(abcdefg_f08_eg0_ab_cdefghijklm[49]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_36_1(abcdefg_f10_eg2_ab_fghijklm[36]),
    .abcd_efgh_ijklmno_f05_out_h_2(abcdefg_f05_a_zxdf[0]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_cc(abcdefg_f09_eg1_ab_cdefghijklm[41]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_3_1(abcdefg_f11_eg3_ab_fghijklm[3]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_ff_1(abcdefg_f11_eg3_ab_a_fghi[8]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_19_2(abcdefg_f11_eg3_ab_fghijklm[19]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_bi_1(abcdefg_f11_eg3_ab_a_fghi[45]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_49_1(abcdefg_f08_eg0_ab_fghijklm[49]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_ee_1(abcdefg_f10_eg2_ab_cdefghijklm[19]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_29_1(abcdefg_f08_eg0_ab_fghijklm[29]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_29_1(abcdefg_f09_eg1_ab_fghijklm[29]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_ed(abcdefg_f09_eg1_ab_cdefghijklm[20]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_de(abcdefg_f09_eg1_ab_cdefghijklm[29]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_dg_2(abcdefg_f10_eg2_ab_a_fghi[27]),
    .abcd_efgh_ijklmno_f04_oilouull_o_2_1(abcdefg_f04_oilouull[2]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_eb_2(abcdefg_f10_eg2_ab_a_fghi[22]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_ea_2(abcdefg_f11_eg3_ab_cdefghijklm[23]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_fc_1(abcdefg_f10_eg2_ab_cdefghijklm[11]),
    .abcd_efgh_ijklmno_f06_out_g(abcdefg_f06_clroilouull[1]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_61_1(abcdefg_f09_eg1_ab_fghijklm[61]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_ee_2(abcdefg_f10_eg2_ab_a_fghi[19]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_47_1(abcdefg_f11_eg3_ab_fghijklm[47]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_36_1(abcdefg_f08_eg0_ab_fghijklm[36]),
    .abcd_efgh_ijklmno_f07_oilouull_o_0_1(abcdefg_f07_oilouull[0]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_j_1(abcdefg_f11_eg3_ab_a_fghi[54]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_52_1(abcdefg_f08_eg0_ab_fghijklm[52]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_gd_1(abcdefg_f11_eg3_ab_a_fghi[0]),
    .abcd_efgh_ijklmno_f07_out_h_2(abcdefg_f07_a_zxdf[0]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_cg_1(abcdefg_f09_eg1_ab_a_fghi[37]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_8_1(abcdefg_f10_eg2_ab_fghijklm[8]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_fh_1(abcdefg_f11_eg3_ab_a_fghi[6]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_52_1(abcdefg_f09_eg1_ab_fghijklm[52]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_ci_2(abcdefg_f11_eg3_ab_cdefghijklm[35]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_15_1(abcdefg_f10_eg2_ab_fghijklm[15]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_df(abcdefg_f09_eg1_ab_cdefghijklm[28]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_ee(abcdefg_f09_eg1_ab_cdefghijklm[19]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_bd_1(abcdefg_f11_eg3_ab_a_fghi[50]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_fe_1(abcdefg_f11_eg3_ab_a_fghi[9]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_di_2(abcdefg_f08_eg0_ab_a_fghi[25]),
    .abcd_efgh_ijklmno_f00_out_d(abcdefg_f00_clroilouull[4]),
    .abcd_efgh_ijklmno_f07_oilouull_o_5_1(abcdefg_f07_oilouull[5]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_41_1(abcdefg_f09_eg1_ab_fghijklm[41]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_cf_2(abcdefg_f08_eg0_ab_cdefghijklm[38]),
    .abcd_efgh_ijklmno_f05_out_b_3(abcdefg_f05_a_zxdf[6]),
    .abcd_efgh_ijklmno_f03_oilouull_o_1_1(abcdefg_f03_oilouull[1]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_dg_1(abcdefg_f09_eg1_ab_a_fghi[27]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_eg(abcdefg_f09_eg1_ab_cdefghijklm[17]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_ce_1(abcdefg_f09_eg1_ab_a_fghi[39]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_fi_2(abcdefg_f11_eg3_ab_cdefghijklm[5]),
    .abcd_efgh_ijklmno_f05_out_g(abcdefg_f05_clroilouull[1]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_bj_2(abcdefg_f10_eg2_ab_cdefghijklm[44]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_db(abcdefg_f09_eg1_ab_cdefghijklm[32]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_g_1(abcdefg_f09_eg1_ab_a_fghi[57]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_bf_2(abcdefg_f08_eg0_ab_cdefghijklm[48]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_bh_2(abcdefg_f08_eg0_ab_cdefghijklm[46]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_23_1(abcdefg_f10_eg2_ab_fghijklm[23]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_61_1(abcdefg_f10_eg2_ab_fghijklm[61]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_db_1(abcdefg_f09_eg1_ab_a_fghi[32]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_f(abcdefg_f09_eg1_ab_cdefghijklm[58]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_57_1(abcdefg_f09_eg1_ab_fghijklm[57]),
    .abcd_efgh_ijklmno_f01_oilouull_o_1_1(abcdefg_f01_oilouull[1]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_eh_2(abcdefg_f08_eg0_ab_a_fghi[16]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_41_1(abcdefg_f11_eg3_ab_fghijklm[41]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_c_2(abcdefg_f08_eg0_ab_cdefghijklm[61]),
    .abcd_efgh_ijklmno_f06_out_e(abcdefg_f06_clroilouull[3]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_ej_1(abcdefg_f11_eg3_ab_a_fghi[14]),
    .abcd_efgh_ijklmno_f02_oilouull_o_1_1(abcdefg_f02_oilouull[1]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_bd_2(abcdefg_f11_eg3_ab_cdefghijklm[50]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_6_1(abcdefg_f08_eg0_ab_fghijklm[6]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_ee_1(abcdefg_f09_eg1_ab_a_fghi[19]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_fc_2(abcdefg_f11_eg3_ab_cdefghijklm[11]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_bd_3(abcdefg_f10_eg2_ab_a_fghi[50]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_df_1(abcdefg_f08_eg0_ab_cdefghijklm[28]),
    .abcd_efgh_ijklmno_f03_out_a(abcdefg_f03_clroilouull[7]),
    .abcd_efgh_ijklmno_f02_oilouull_o_0_1(abcdefg_f02_oilouull[0]),
    .abcd_efgh_ijklmno_f00_out_g_2(abcdefg_f00_a_zxdf[1]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_43_1(abcdefg_f08_eg0_ab_fghijklm[43]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_59_1(abcdefg_f08_eg0_ab_fghijklm[59]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_ff_1(abcdefg_f09_eg1_ab_a_fghi[8]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_bh_2(abcdefg_f10_eg2_ab_cdefghijklm[46]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_0_1(abcdefg_f09_eg1_ab_fghijklm[0]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_ec_2(abcdefg_f08_eg0_ab_a_fghi[21]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_33_1(abcdefg_f09_eg1_ab_fghijklm[33]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_fh_1(abcdefg_f09_eg1_ab_a_fghi[6]),
    .abcd_efgh_ijklmno_f02_oilouull_o_4_1(abcdefg_f02_oilouull[4]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_31_1(abcdefg_f10_eg2_ab_fghijklm[31]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_fa_1(abcdefg_f10_eg2_ab_cdefghijklm[13]),
    .abcd_efgh_ijklmno_f05_out_f(abcdefg_f05_clroilouull[2]),
    .abcd_efgh_ijklmno_f04_out_e_2(abcdefg_f04_a_zxdf[3]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_dd_1(abcdefg_f09_eg1_ab_a_fghi[30]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_12_1(abcdefg_f11_eg3_ab_fghijklm[12]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_bf_1(abcdefg_f09_eg1_ab_a_fghi[48]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_23_1(abcdefg_f08_eg0_ab_fghijklm[23]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_dj_2(abcdefg_f08_eg0_ab_a_fghi[24]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_ci_3(abcdefg_f10_eg2_ab_a_fghi[35]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_17_1(abcdefg_f08_eg0_ab_fghijklm[17]),
    .abcd_efgh_ijklmno_f02_out_f_2(abcdefg_f02_a_zxdf[2]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_bb_1(abcdefg_f11_eg3_ab_a_fghi[52]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_cc_1(abcdefg_f11_eg3_ab_a_fghi[41]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_f_1(abcdefg_f11_eg3_ab_a_fghi[58]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_fi(abcdefg_f09_eg1_ab_cdefghijklm[5]),
    .abcd_efgh_ijklmno_f03_out_h(abcdefg_f03_clroilouull[0]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_e_1(abcdefg_f11_eg3_ab_a_fghi[59]),
    .abcd_efgh_ijklmno_f01_out_b_3(abcdefg_f01_a_zxdf[6]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_55_1(abcdefg_f08_eg0_ab_fghijklm[55]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_bj_3(abcdefg_f10_eg2_ab_a_fghi[44]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_d_2(abcdefg_f08_eg0_ab_cdefghijklm[60]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_bi_3(abcdefg_f08_eg0_ab_a_fghi[45]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_fg_1(abcdefg_f09_eg1_ab_a_fghi[7]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_ej_2(abcdefg_f10_eg2_ab_a_fghi[14]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_cb_2(abcdefg_f08_eg0_ab_cdefghijklm[42]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_fi_1(abcdefg_f10_eg2_ab_cdefghijklm[5]),
    .abcd_efgh_ijklmno_f01_out_c(abcdefg_f01_clroilouull[5]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_fa_2(abcdefg_f11_eg3_ab_cdefghijklm[13]),
    .abcd_efgh_ijklmno_f07_out_b_3(abcdefg_f07_a_zxdf[6]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_2_1(abcdefg_f09_eg1_ab_fghijklm[2]),
    .abcd_efgh_ijklmno_f07_oilouull_o_2_1(abcdefg_f07_oilouull[2]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_ed_2(abcdefg_f10_eg2_ab_a_fghi[20]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_32_1(abcdefg_f08_eg0_ab_fghijklm[32]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_29_1(abcdefg_f10_eg2_ab_fghijklm[29]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_ef_1(abcdefg_f11_eg3_ab_a_fghi[18]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_15_1(abcdefg_f09_eg1_ab_fghijklm[15]),
    .abcd_efgh_ijklmno_f04_out_c_2(abcdefg_f04_a_zxdf[5]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_cd(abcdefg_f09_eg1_ab_cdefghijklm[40]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_57_1(abcdefg_f08_eg0_ab_fghijklm[57]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_ee_2(abcdefg_f11_eg3_ab_cdefghijklm[19]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_3_1(abcdefg_f09_eg1_ab_fghijklm[3]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_20_1(abcdefg_f10_eg2_ab_fghijklm[20]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_16_1(abcdefg_f08_eg0_ab_fghijklm[16]),
    .abcd_efgh_ijklmno_f06_oilouull_o_1_1(abcdefg_f06_oilouull[1]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_cg(abcdefg_f09_eg1_ab_cdefghijklm[37]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_cd_3(abcdefg_f10_eg2_ab_a_fghi[40]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_35_1(abcdefg_f10_eg2_ab_fghijklm[35]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_j_3(abcdefg_f10_eg2_ab_a_fghi[54]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_dc_2(abcdefg_f10_eg2_ab_a_fghi[31]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_34_1(abcdefg_f08_eg0_ab_fghijklm[34]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_bi_2(abcdefg_f10_eg2_ab_cdefghijklm[45]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_48_1(abcdefg_f09_eg1_ab_fghijklm[48]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_1_2(abcdefg_f10_eg2_ab_fghijklm[1]),
    .abcd_efgh_ijklmno_f07_out_g(abcdefg_f07_clroilouull[1]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_c_2(abcdefg_f11_eg3_ab_cdefghijklm[61]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_24_1(abcdefg_f10_eg2_ab_fghijklm[24]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_fj_2(abcdefg_f10_eg2_ab_a_fghi[4]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_bi_1(abcdefg_f09_eg1_ab_a_fghi[45]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_eb_2(abcdefg_f11_eg3_ab_cdefghijklm[22]),
    .abcd_efgh_ijklmno_f00_oilouull_o_5_1(abcdefg_f00_oilouull[5]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_30_1(abcdefg_f08_eg0_ab_fghijklm[30]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_11_1(abcdefg_f11_eg3_ab_fghijklm[11]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_26_1(abcdefg_f11_eg3_ab_fghijklm[26]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_45_1(abcdefg_f08_eg0_ab_fghijklm[45]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_dj_1(abcdefg_f10_eg2_ab_cdefghijklm[24]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_gd_1(abcdefg_f10_eg2_ab_cdefghijklm[0]),
    .abcd_efgh_ijklmno_f05_out_b(abcdefg_f05_clroilouull[6]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_ef_2(abcdefg_f08_eg0_ab_a_fghi[18]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_dg(abcdefg_f09_eg1_ab_cdefghijklm[27]),
    .abcd_efgh_ijklmno_f02_oilouull_o_6_2(abcdefg_f02_oilouull[6]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_39_1(abcdefg_f11_eg3_ab_fghijklm[39]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_bh_3(abcdefg_f10_eg2_ab_a_fghi[46]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_fc_1(abcdefg_f08_eg0_ab_cdefghijklm[11]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_fa(abcdefg_f09_eg1_ab_cdefghijklm[13]),
    .abcd_efgh_ijklmno_f04_out_b_3(abcdefg_f04_a_zxdf[6]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_21_1(abcdefg_f08_eg0_ab_fghijklm[21]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_bc_3(abcdefg_f08_eg0_ab_a_fghi[51]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_dd_1(abcdefg_f08_eg0_ab_cdefghijklm[30]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_fc_1(abcdefg_f09_eg1_ab_a_fghi[11]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_22_1(abcdefg_f11_eg3_ab_fghijklm[22]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_14_1(abcdefg_f11_eg3_ab_fghijklm[14]),
    .abcd_efgh_ijklmno_f02_out_d_2(abcdefg_f02_a_zxdf[4]),
    .abcd_efgh_ijklmno_f06_out_h(abcdefg_f06_clroilouull[0]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_37_1(abcdefg_f09_eg1_ab_fghijklm[37]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_eh_1(abcdefg_f09_eg1_ab_a_fghi[16]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_12_1(abcdefg_f09_eg1_ab_fghijklm[12]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_cd_1(abcdefg_f09_eg1_ab_a_fghi[40]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_60_1(abcdefg_f11_eg3_ab_fghijklm[60]),
    .abcd_efgh_ijklmno_f03_out_f_2(abcdefg_f03_a_zxdf[2]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_43_1(abcdefg_f11_eg3_ab_fghijklm[43]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_dc_2(abcdefg_f08_eg0_ab_a_fghi[31]),
    .abcd_efgh_ijklmno_f07_out_b(abcdefg_f07_clroilouull[6]),
    .abcd_efgh_ijklmno_f03_out_b_3(abcdefg_f03_a_zxdf[6]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_ea_1(abcdefg_f10_eg2_ab_cdefghijklm[23]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_eg_1(abcdefg_f08_eg0_ab_cdefghijklm[17]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_fc_2(abcdefg_f08_eg0_ab_a_fghi[11]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_gc_1(abcdefg_f08_eg0_ab_cdefghijklm[1]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_da(abcdefg_f09_eg1_ab_cdefghijklm[33]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_gb_2(abcdefg_f11_eg3_ab_cdefghijklm[2]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_ba_2(abcdefg_f10_eg2_ab_cdefghijklm[53]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_fb_2(abcdefg_f10_eg2_ab_a_fghi[12]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_ee_1(abcdefg_f11_eg3_ab_a_fghi[19]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_32_1(abcdefg_f09_eg1_ab_fghijklm[32]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_gc_2(abcdefg_f11_eg3_ab_cdefghijklm[1]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_ee_1(abcdefg_f08_eg0_ab_cdefghijklm[19]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_36_1(abcdefg_f09_eg1_ab_fghijklm[36]),
    .abcd_efgh_ijklmno_f02_out_a(abcdefg_f02_clroilouull[7]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_9_1(abcdefg_f08_eg0_ab_fghijklm[9]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_5_1(abcdefg_f09_eg1_ab_fghijklm[5]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_bh_2(abcdefg_f11_eg3_ab_cdefghijklm[46]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_35_1(abcdefg_f09_eg1_ab_fghijklm[35]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_ca(abcdefg_f09_eg1_ab_cdefghijklm[43]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_47_1(abcdefg_f08_eg0_ab_fghijklm[47]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_gc_1(abcdefg_f11_eg3_ab_a_fghi[1]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_ba_2(abcdefg_f08_eg0_ab_cdefghijklm[53]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_44_1(abcdefg_f11_eg3_ab_fghijklm[44]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_9_1(abcdefg_f09_eg1_ab_fghijklm[9]),
    .abcd_efgh_ijklmno_f00_oilouull_o_3_1(abcdefg_f00_oilouull[3]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_fe_2(abcdefg_f11_eg3_ab_cdefghijklm[9]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_ec_1(abcdefg_f09_eg1_ab_a_fghi[21]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_de_2(abcdefg_f10_eg2_ab_a_fghi[29]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_29_1(abcdefg_f11_eg3_ab_fghijklm[29]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_g_3(abcdefg_f08_eg0_ab_a_fghi[57]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_fi_2(abcdefg_f10_eg2_ab_a_fghi[5]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_27_1(abcdefg_f08_eg0_ab_fghijklm[27]),
    .abcd_efgh_ijklmno_f11_eg3_ge_out_fc_1(abcdefg_f11_eg3_ab_a_fghi[11]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_42_1(abcdefg_f10_eg2_ab_fghijklm[42]),
    .abcd_efgh_ijklmno_f04_oilouull_o_4_1(abcdefg_f04_oilouull[4]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_30_1(abcdefg_f09_eg1_ab_fghijklm[30]),
    .abcd_efgh_ijklmno_f01_oilouull_o_3_1(abcdefg_f01_oilouull[3]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_fj_1(abcdefg_f10_eg2_ab_cdefghijklm[4]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_55_1(abcdefg_f11_eg3_ab_fghijklm[55]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_42_1(abcdefg_f08_eg0_ab_fghijklm[42]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_gd(abcdefg_f09_eg1_ab_cdefghijklm[0]),
    .abcd_efgh_ijklmno_f09_eg1_ge_out_eg_1(abcdefg_f09_eg1_ab_a_fghi[17]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_8_1(abcdefg_f08_eg0_ab_fghijklm[8]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_50_1(abcdefg_f11_eg3_ab_fghijklm[50]),
    .abcd_efgh_ijklmno_f06_out_f_2(abcdefg_f06_a_zxdf[2]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_26_1(abcdefg_f09_eg1_ab_fghijklm[26]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_30_1(abcdefg_f11_eg3_ab_fghijklm[30]),
    .abcd_efgh_ijklmno_f10_eg2_ab_fghijklm_o_55_1(abcdefg_f10_eg2_ab_fghijklm[55]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_df_2(abcdefg_f08_eg0_ab_a_fghi[28]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_28_1(abcdefg_f09_eg1_ab_fghijklm[28]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_22_1(abcdefg_f09_eg1_ab_fghijklm[22]),
    .abcd_efgh_ijklmno_f09_eg1_ab_fghijklm_o_45_1(abcdefg_f09_eg1_ab_fghijklm[45]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_46_1(abcdefg_f08_eg0_ab_fghijklm[46]),
    .abcd_efgh_ijklmno_f01_out_f(abcdefg_f01_clroilouull[2]),
    .abcd_efgh_ijklmno_f11_eg3_ab_fghijklm_o_36_1(abcdefg_f11_eg3_ab_fghijklm[36]),
    .abcd_efgh_ijklmno_f05_out_f_2(abcdefg_f05_a_zxdf[2]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_ch_2(abcdefg_f08_eg0_ab_cdefghijklm[36]),
    .abcd_efgh_ijklmno_f10_eg2_ge_out_cj_3(abcdefg_f10_eg2_ab_a_fghi[34]),
    .abcd_efgh_ijklmno_f04_oilouull_o_3_1(abcdefg_f04_oilouull[3]),
    .abcd_efgh_ijklmno_f08_eg0_ge_out_cd_3(abcdefg_f08_eg0_ab_a_fghi[40]),
    .abcd_efgh_ijklmno_f08_eg0_ab_fghijklm_o_56_1(abcdefg_f08_eg0_ab_fghijklm[56]),
    
    
    );*/
   TEST TEST (/*AUTOINST*/);
   
endmodule

module TEST (/*AUTOARG*/);
   parameter NO = 6456;
endmodule
