module foo;
   modport foo_mp;
   modport foo_mp1(a);
   modport foo_mp2(clocking bar_cb);
   a;
endmodule // foo
