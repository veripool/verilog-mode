// msg2404

module top
  (
   /*AUTOINPUT*/
   /*AUTOOUTPUT*/
   );

   /*AUTOLOGIC*/

   submod inst
     (/*AUTOINST*/);
    
endmodule

module submod
  (input [2*2:1] x);
endmodule

// Local Variables:
// verilog-auto-simplify-expressions: nil
// End:
