
module flag_f_reeves
  (/*AUTOARG*/) ;

   /*AUTOOUTPUT*/

   /*AUTOINPUT*/

   flag_f_reeves_IBUF ibuf
     (/*AUTOINST*/);

endmodule
// Local Variables:
// verilog-library-flags: ("-F subdir/flag_frel_reeves.vc")
// End:
