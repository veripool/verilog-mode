`include "x.h"
//
module x;
   ////
   reg             y;
endmodule // x
