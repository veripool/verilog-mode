module flag_f_reeves_IBUF (input a, output q);
endmodule
