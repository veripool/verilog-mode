module autoinoutin (/*AUTOARG*/);

   /*AUTOINOUTIN("inst")*/

endmodule

