module indent_enum;
   
   enum int unsigned {
      STATE_0 = 0,
      STATE_2 = 2
   } state;
   
   enum int unsigned {
      STATE_0 = 0,
      STATE_1,
      STATE_2
   } state, next;
   
endmodule
