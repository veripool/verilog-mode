// issue 1080 - Indentation of a virtual class definition after a typedef class line
typedef class foo;
virtual class bar;
endclass : bar
